// Computer_System_D5M_Subsystem.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module Computer_System_D5M_Subsystem (
		input  wire [1:0]  avalon_d5m_config_slave_address,       //    avalon_d5m_config_slave.address
		input  wire [3:0]  avalon_d5m_config_slave_byteenable,    //                           .byteenable
		input  wire        avalon_d5m_config_slave_read,          //                           .read
		input  wire        avalon_d5m_config_slave_write,         //                           .write
		input  wire [31:0] avalon_d5m_config_slave_writedata,     //                           .writedata
		output wire [31:0] avalon_d5m_config_slave_readdata,      //                           .readdata
		output wire        avalon_d5m_config_slave_waitrequest,   //                           .waitrequest
		inout  wire        d5m_config_I2C_SDAT,                   //                 d5m_config.I2C_SDAT
		output wire        d5m_config_I2C_SCLK,                   //                           .I2C_SCLK
		input  wire [15:0] d5m_config_exposure,                   //                           .exposure
		input  wire        sys_clk_clk,                           //                    sys_clk.clk
		input  wire        sys_reset_reset_n,                     //                  sys_reset.reset_n
		input  wire        video_in_PIXEL_CLK,                    //                   video_in.PIXEL_CLK
		input  wire        video_in_LINE_VALID,                   //                           .LINE_VALID
		input  wire        video_in_FRAME_VALID,                  //                           .FRAME_VALID
		input  wire        video_in_pixel_clk_reset,              //                           .pixel_clk_reset
		input  wire [11:0] video_in_PIXEL_DATA,                   //                           .PIXEL_DATA
		input  wire [1:0]  video_in_dma_control_slave_address,    // video_in_dma_control_slave.address
		input  wire [3:0]  video_in_dma_control_slave_byteenable, //                           .byteenable
		input  wire        video_in_dma_control_slave_read,       //                           .read
		input  wire        video_in_dma_control_slave_write,      //                           .write
		input  wire [31:0] video_in_dma_control_slave_writedata,  //                           .writedata
		output wire [31:0] video_in_dma_control_slave_readdata,   //                           .readdata
		output wire [31:0] video_in_dma_master_address,           //        video_in_dma_master.address
		input  wire        video_in_dma_master_waitrequest,       //                           .waitrequest
		output wire        video_in_dma_master_write,             //                           .write
		output wire [15:0] video_in_dma_master_writedata          //                           .writedata
	);

	wire         bayer_resampler_avalon_bayer_source_valid;              // Bayer_Resampler:stream_out_valid -> Video_In_RGB_Resampler:stream_in_valid
	wire  [23:0] bayer_resampler_avalon_bayer_source_data;               // Bayer_Resampler:stream_out_data -> Video_In_RGB_Resampler:stream_in_data
	wire         bayer_resampler_avalon_bayer_source_ready;              // Video_In_RGB_Resampler:stream_in_ready -> Bayer_Resampler:stream_out_ready
	wire         bayer_resampler_avalon_bayer_source_startofpacket;      // Bayer_Resampler:stream_out_startofpacket -> Video_In_RGB_Resampler:stream_in_startofpacket
	wire         bayer_resampler_avalon_bayer_source_endofpacket;        // Bayer_Resampler:stream_out_endofpacket -> Video_In_RGB_Resampler:stream_in_endofpacket
	wire         video_in_clipper_avalon_clipper_source_valid;           // Video_In_Clipper:stream_out_valid -> Video_In_Scaler:stream_in_valid
	wire  [15:0] video_in_clipper_avalon_clipper_source_data;            // Video_In_Clipper:stream_out_data -> Video_In_Scaler:stream_in_data
	wire         video_in_clipper_avalon_clipper_source_ready;           // Video_In_Scaler:stream_in_ready -> Video_In_Clipper:stream_out_ready
	wire         video_in_clipper_avalon_clipper_source_startofpacket;   // Video_In_Clipper:stream_out_startofpacket -> Video_In_Scaler:stream_in_startofpacket
	wire         video_in_clipper_avalon_clipper_source_endofpacket;     // Video_In_Clipper:stream_out_endofpacket -> Video_In_Scaler:stream_in_endofpacket
	wire         video_in_avalon_decoder_source_valid;                   // Video_In:stream_out_valid -> Bayer_Resampler:stream_in_valid
	wire   [7:0] video_in_avalon_decoder_source_data;                    // Video_In:stream_out_data -> Bayer_Resampler:stream_in_data
	wire         video_in_avalon_decoder_source_ready;                   // Bayer_Resampler:stream_in_ready -> Video_In:stream_out_ready
	wire         video_in_avalon_decoder_source_startofpacket;           // Video_In:stream_out_startofpacket -> Bayer_Resampler:stream_in_startofpacket
	wire         video_in_avalon_decoder_source_endofpacket;             // Video_In:stream_out_endofpacket -> Bayer_Resampler:stream_in_endofpacket
	wire         video_in_rgb_resampler_avalon_rgb_source_valid;         // Video_In_RGB_Resampler:stream_out_valid -> Video_In_Clipper:stream_in_valid
	wire  [15:0] video_in_rgb_resampler_avalon_rgb_source_data;          // Video_In_RGB_Resampler:stream_out_data -> Video_In_Clipper:stream_in_data
	wire         video_in_rgb_resampler_avalon_rgb_source_ready;         // Video_In_Clipper:stream_in_ready -> Video_In_RGB_Resampler:stream_out_ready
	wire         video_in_rgb_resampler_avalon_rgb_source_startofpacket; // Video_In_RGB_Resampler:stream_out_startofpacket -> Video_In_Clipper:stream_in_startofpacket
	wire         video_in_rgb_resampler_avalon_rgb_source_endofpacket;   // Video_In_RGB_Resampler:stream_out_endofpacket -> Video_In_Clipper:stream_in_endofpacket
	wire         video_in_scaler_avalon_scaler_source_valid;             // Video_In_Scaler:stream_out_valid -> Video_In_DMA:stream_valid
	wire  [15:0] video_in_scaler_avalon_scaler_source_data;              // Video_In_Scaler:stream_out_data -> Video_In_DMA:stream_data
	wire         video_in_scaler_avalon_scaler_source_ready;             // Video_In_DMA:stream_ready -> Video_In_Scaler:stream_out_ready
	wire         video_in_scaler_avalon_scaler_source_startofpacket;     // Video_In_Scaler:stream_out_startofpacket -> Video_In_DMA:stream_startofpacket
	wire         video_in_scaler_avalon_scaler_source_endofpacket;       // Video_In_Scaler:stream_out_endofpacket -> Video_In_DMA:stream_endofpacket
	wire         rst_controller_reset_out_reset;                         // rst_controller:reset_out -> [Bayer_Resampler:reset, D5M_Config:reset, Video_In:reset, Video_In_Clipper:reset, Video_In_DMA:reset, Video_In_RGB_Resampler:reset, Video_In_Scaler:reset]

	Computer_System_D5M_Subsystem_Bayer_Resampler bayer_resampler (
		.clk                      (sys_clk_clk),                                       //                 clk.clk
		.reset                    (rst_controller_reset_out_reset),                    //               reset.reset
		.stream_in_data           (video_in_avalon_decoder_source_data),               //   avalon_bayer_sink.data
		.stream_in_startofpacket  (video_in_avalon_decoder_source_startofpacket),      //                    .startofpacket
		.stream_in_endofpacket    (video_in_avalon_decoder_source_endofpacket),        //                    .endofpacket
		.stream_in_valid          (video_in_avalon_decoder_source_valid),              //                    .valid
		.stream_in_ready          (video_in_avalon_decoder_source_ready),              //                    .ready
		.stream_out_ready         (bayer_resampler_avalon_bayer_source_ready),         // avalon_bayer_source.ready
		.stream_out_data          (bayer_resampler_avalon_bayer_source_data),          //                    .data
		.stream_out_startofpacket (bayer_resampler_avalon_bayer_source_startofpacket), //                    .startofpacket
		.stream_out_endofpacket   (bayer_resampler_avalon_bayer_source_endofpacket),   //                    .endofpacket
		.stream_out_valid         (bayer_resampler_avalon_bayer_source_valid)          //                    .valid
	);

	Computer_System_D5M_Subsystem_D5M_Config d5m_config (
		.clk         (sys_clk_clk),                         //                    clk.clk
		.reset       (rst_controller_reset_out_reset),      //                  reset.reset
		.address     (avalon_d5m_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (avalon_d5m_config_slave_byteenable),  //                       .byteenable
		.read        (avalon_d5m_config_slave_read),        //                       .read
		.write       (avalon_d5m_config_slave_write),       //                       .write
		.writedata   (avalon_d5m_config_slave_writedata),   //                       .writedata
		.readdata    (avalon_d5m_config_slave_readdata),    //                       .readdata
		.waitrequest (avalon_d5m_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (d5m_config_I2C_SDAT),                 //     external_interface.export
		.I2C_SCLK    (d5m_config_I2C_SCLK),                 //                       .export
		.exposure    (d5m_config_exposure)                  //                       .export
	);

	Computer_System_D5M_Subsystem_Video_In video_in (
		.clk                      (sys_clk_clk),                                  //                   clk.clk
		.reset                    (rst_controller_reset_out_reset),               //                 reset.reset
		.stream_out_ready         (video_in_avalon_decoder_source_ready),         // avalon_decoder_source.ready
		.stream_out_startofpacket (video_in_avalon_decoder_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (video_in_avalon_decoder_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (video_in_avalon_decoder_source_valid),         //                      .valid
		.stream_out_data          (video_in_avalon_decoder_source_data),          //                      .data
		.PIXEL_CLK                (video_in_PIXEL_CLK),                           //    external_interface.export
		.LINE_VALID               (video_in_LINE_VALID),                          //                      .export
		.FRAME_VALID              (video_in_FRAME_VALID),                         //                      .export
		.pixel_clk_reset          (video_in_pixel_clk_reset),                     //                      .export
		.PIXEL_DATA               (video_in_PIXEL_DATA)                           //                      .export
	);

	Computer_System_D5M_Subsystem_Video_In_Clipper video_in_clipper (
		.clk                      (sys_clk_clk),                                            //                   clk.clk
		.reset                    (rst_controller_reset_out_reset),                         //                 reset.reset
		.stream_in_data           (video_in_rgb_resampler_avalon_rgb_source_data),          //   avalon_clipper_sink.data
		.stream_in_startofpacket  (video_in_rgb_resampler_avalon_rgb_source_startofpacket), //                      .startofpacket
		.stream_in_endofpacket    (video_in_rgb_resampler_avalon_rgb_source_endofpacket),   //                      .endofpacket
		.stream_in_valid          (video_in_rgb_resampler_avalon_rgb_source_valid),         //                      .valid
		.stream_in_ready          (video_in_rgb_resampler_avalon_rgb_source_ready),         //                      .ready
		.stream_out_ready         (video_in_clipper_avalon_clipper_source_ready),           // avalon_clipper_source.ready
		.stream_out_data          (video_in_clipper_avalon_clipper_source_data),            //                      .data
		.stream_out_startofpacket (video_in_clipper_avalon_clipper_source_startofpacket),   //                      .startofpacket
		.stream_out_endofpacket   (video_in_clipper_avalon_clipper_source_endofpacket),     //                      .endofpacket
		.stream_out_valid         (video_in_clipper_avalon_clipper_source_valid)            //                      .valid
	);

	Computer_System_D5M_Subsystem_Video_In_DMA video_in_dma (
		.clk                  (sys_clk_clk),                                        //                      clk.clk
		.reset                (rst_controller_reset_out_reset),                     //                    reset.reset
		.stream_data          (video_in_scaler_avalon_scaler_source_data),          //          avalon_dma_sink.data
		.stream_startofpacket (video_in_scaler_avalon_scaler_source_startofpacket), //                         .startofpacket
		.stream_endofpacket   (video_in_scaler_avalon_scaler_source_endofpacket),   //                         .endofpacket
		.stream_valid         (video_in_scaler_avalon_scaler_source_valid),         //                         .valid
		.stream_ready         (video_in_scaler_avalon_scaler_source_ready),         //                         .ready
		.slave_address        (video_in_dma_control_slave_address),                 // avalon_dma_control_slave.address
		.slave_byteenable     (video_in_dma_control_slave_byteenable),              //                         .byteenable
		.slave_read           (video_in_dma_control_slave_read),                    //                         .read
		.slave_write          (video_in_dma_control_slave_write),                   //                         .write
		.slave_writedata      (video_in_dma_control_slave_writedata),               //                         .writedata
		.slave_readdata       (video_in_dma_control_slave_readdata),                //                         .readdata
		.master_address       (video_in_dma_master_address),                        //        avalon_dma_master.address
		.master_waitrequest   (video_in_dma_master_waitrequest),                    //                         .waitrequest
		.master_write         (video_in_dma_master_write),                          //                         .write
		.master_writedata     (video_in_dma_master_writedata)                       //                         .writedata
	);

	Computer_System_D5M_Subsystem_Video_In_RGB_Resampler video_in_rgb_resampler (
		.clk                      (sys_clk_clk),                                            //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                         //             reset.reset
		.stream_in_startofpacket  (bayer_resampler_avalon_bayer_source_startofpacket),      //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (bayer_resampler_avalon_bayer_source_endofpacket),        //                  .endofpacket
		.stream_in_valid          (bayer_resampler_avalon_bayer_source_valid),              //                  .valid
		.stream_in_ready          (bayer_resampler_avalon_bayer_source_ready),              //                  .ready
		.stream_in_data           (bayer_resampler_avalon_bayer_source_data),               //                  .data
		.stream_out_ready         (video_in_rgb_resampler_avalon_rgb_source_ready),         // avalon_rgb_source.ready
		.stream_out_startofpacket (video_in_rgb_resampler_avalon_rgb_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (video_in_rgb_resampler_avalon_rgb_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (video_in_rgb_resampler_avalon_rgb_source_valid),         //                  .valid
		.stream_out_data          (video_in_rgb_resampler_avalon_rgb_source_data)           //                  .data
	);

	Computer_System_D5M_Subsystem_Video_In_Scaler video_in_scaler (
		.clk                      (sys_clk_clk),                                          //                  clk.clk
		.reset                    (rst_controller_reset_out_reset),                       //                reset.reset
		.stream_in_startofpacket  (video_in_clipper_avalon_clipper_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (video_in_clipper_avalon_clipper_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (video_in_clipper_avalon_clipper_source_valid),         //                     .valid
		.stream_in_ready          (video_in_clipper_avalon_clipper_source_ready),         //                     .ready
		.stream_in_data           (video_in_clipper_avalon_clipper_source_data),          //                     .data
		.stream_out_ready         (video_in_scaler_avalon_scaler_source_ready),           // avalon_scaler_source.ready
		.stream_out_startofpacket (video_in_scaler_avalon_scaler_source_startofpacket),   //                     .startofpacket
		.stream_out_endofpacket   (video_in_scaler_avalon_scaler_source_endofpacket),     //                     .endofpacket
		.stream_out_valid         (video_in_scaler_avalon_scaler_source_valid),           //                     .valid
		.stream_out_data          (video_in_scaler_avalon_scaler_source_data)             //                     .data
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~sys_reset_reset_n),             // reset_in0.reset
		.clk            (sys_clk_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
